module BCD (input [3:0] BINARY,
				output reg [6:0] SEGMENTS);
				
always@(*)
	case(BINARY)
		0:SEGMENTS=7'b1000000;
		1:SEGMENTS=7'b1111001;
		2:SEGMENTS=7'b0100100;
		3:SEGMENTS=7'b0110000;
		4:SEGMENTS=7'b0011001;
		5:SEGMENTS=7'b0010010;
		6:SEGMENTS=7'b0000010;
		7:SEGMENTS=7'b1111000;
		8:SEGMENTS=7'b0000000;
		9:SEGMENTS=7'b0010000;
		10:SEGMENTS=7'b0001000;
		11:SEGMENTS=7'b0000011;
		12:SEGMENTS=7'b1000110;
		13:SEGMENTS=7'b0100001;
		14:SEGMENTS=7'b0000110;
		15:SEGMENTS=7'b0001110;
		default:SEGMENTS=7'b1111111;
	endcase
	
endmodule 