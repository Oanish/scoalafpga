module top(
    input wire CLK,             // board clock: 100 MHz on Arty & Basys 3
    input wire RST_BTN,         // reset button
    output wire VGA_HS_O,       // horizontal sync output
    output wire VGA_VS_O,       // vertical sync output
    output wire [3:0] VGA_R,    // 4-bit VGA red output
    output wire [3:0] VGA_G,    // 4-bit VGA green output
    output wire [3:0] VGA_B     // 4-bit VGA blue output
    );

    wire rst = ~RST_BTN;  // reset is active low on Arty

    // generate a 25 MHz pixel strobe
    reg [15:0] cnt;
    reg pix_stb;
    always @(posedge CLK)
        {pix_stb, cnt} <= cnt + 16'h8000;  // divide by 2: (2^16)/2 = 0x8000

    wire [9:0] x;  // current pixel x position: 10-bit value: 0-1023
    wire [8:0] y;  // current pixel y position:  9-bit value: 0-511

    vga640x480 display (
        .i_clk(CLK),
        .i_pix_stb(pix_stb),
        .i_rst(rst),
        .o_hs(VGA_HS_O), 
        .o_vs(VGA_VS_O), 
        .o_x(x), 
        .o_y(y)
    );

    // Four overlapping squares
    wire sq_a, sq_b, sq_c, sq_d;
    assign sq_a = ((x > 260/*120*/) & (y > 40) & (x < 380/*280*/) & (y < 440/*200*/)) ? 1 : 0;
    assign sq_b = ((x > 120/*260*/) & (y > 180) & (x < 520/*380*/) & (y < 300/*280*/)) ? 1 : 0;
    //assign sq_c = ((x > 280) & (y > 200) & (x < 440) & (y < 360)) ? 1 : 0;
    //assign sq_d = ((x > 360) & (y > 280) & (x < 520) & (y < 440)) ? 1 : 0;

    assign VGA_R = {sq_a | sq_b, sq_a | sq_b, sq_a | sq_b, sq_a | sq_b};//sq_b;         // square b is red
    assign VGA_G = {sq_a | sq_b, 1'b0, 1'b0, 1'b0};  // squares a and d are green
    assign VGA_B = {sq_a | sq_b, 1'b0, sq_a | sq_b, sq_a | sq_b};         // square c is blue
endmodule